`timescale 1ns/10ps
`define SDFFILE     "../02_SYN/Netlist/IOTDF_syn.sdf"     //Modify your sdf file name
`define CYCLE       6.5                   //Modify your CYCLE 
`define DEL         1.0
`define PAT_NUM     64
`define End_CYCLE   1000000 
`define DES_DEBUG


module test;
reg           clk;
reg           rst;
reg           in_en;
reg  [7:0]    iot_in;
reg  [2:0]    fn_sel;
wire          busy;
wire          valid;
wire [127:0]  iot_out;
integer cycle_count;

`ifdef p1
   localparam PAT_NUM = 64;
   localparam F1_NUM = 64;
   localparam F2_NUM = 64;
   localparam F3_NUM = 64;
   localparam F4_NUM = 64;
`elsif p2 // modify the following number according to your pattern
   localparam PAT_NUM = 64;
   localparam F1_NUM = 64;
   localparam F2_NUM = 64;
   localparam F3_NUM = 64;
   localparam F4_NUM = 64;
`else
   localparam PAT_NUM = 64;
   localparam F1_NUM = 64;
   localparam F2_NUM = 64;
   localparam F3_NUM = 64;
   localparam F4_NUM = 64;
`endif


reg  [127:0]  pat_mem[0:PAT_NUM-1];
reg  [127:0]  f1_mem [0:F1_NUM-1];
reg  [127:0]  f2_mem [0:F2_NUM-1];
reg  [127:0]  f3_mem [0:F3_NUM-1];
reg  [127:0]  f4_mem [0:F4_NUM-1];
reg  [127:0]  in_tmp;
reg  [127:0]  out_tmp;
integer       i, j, x, in_l, out_h, out_l, pass, err, err_a;
reg           over, over1, over2;
reg [8*40-1:0] pattern_file_path;
reg [8*34-1:0] func_ans_path;

//wire [3:0] r_load_cnt;
//wire r_state;



IOTDF u_IOTDF( .clk        (clk        ),
               .rst        (rst        ),
               .in_en      (in_en      ), 
               .iot_in     (iot_in     ),
               .fn_sel     (fn_sel     ),
               .busy       (busy       ), 
               .valid      (valid      ), 
               .iot_out    (iot_out    )
               //.r_load_cnt (r_load_cnt),
               //.r_state    (r_state)
             );

/*
`ifdef F4    
               .low        (128'h6FFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF),
               .high       (128'hAFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF),
`elsif F5    
               .low        (128'h7FFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF),
               .high       (128'hBFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF),
`endif
*/

// des debug %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
// `ifdef DES_DEBUG
// // 把 des_core 裡一些重要的訊號拉出來看
// // 注意：這些都是 hierarchical reference，不會影響合成，只用在模擬
// wire [1:0]  des_state    = u_IOTDF.u_des_core.state;
// wire [3:0]  des_round    = u_IOTDF.u_des_core.round_idx;
// wire [31:0] des_L        = u_IOTDF.u_des_core.L_reg;
// wire [31:0] des_R        = u_IOTDF.u_des_core.R_reg;
// wire [31:0] des_f        = u_IOTDF.u_des_core.f_out;
// wire [47:0] des_curkey   = u_IOTDF.u_des_core.cur_subkey;
// wire [63:0] des_ip_out   = u_IOTDF.u_des_core.ip_out;
// wire [55:0] des_pc1_out  = u_IOTDF.u_des_core.pc1_out;
// wire [63:0] des_text_in  = u_IOTDF.u_des_core.text_in;

// // optional: 看 subkey[0] ~ subkey[3] 生成是否正確
// wire [47:0] des_k0 = u_IOTDF.u_des_core.subkey[0];
// wire [47:0] des_k1 = u_IOTDF.u_des_core.subkey[1];
// wire [47:0] des_k2 = u_IOTDF.u_des_core.subkey[2];
// wire [47:0] des_k3 = u_IOTDF.u_des_core.subkey[3];

// // 在 S_KEY 階段，每一輪把 subkey dump 出來
// always @(posedge clk) begin
//     // 只在 F1 (fn_sel=1) 且第一筆 pattern (x==0) 時印，避免太爆
//     if (fn_sel == 3'd1 && x == 0 && des_state == 2'd1) begin
//         $display("[DES KEY] t=%0t round=%2d C=%07h D=%07h subkey=%012h",
//                  $time, des_round, u_IOTDF.u_des_core.C, u_IOTDF.u_des_core.D,
//                  des_curkey);
//     end
// end

// // 在 S_ROUND 階段，每一輪印 L/R + f_out + subkey
// always @(posedge clk) begin
//     if (fn_sel == 3'd1 && x == 0 && des_state == 2'd2) begin
//         $display("[DES ROUND] t=%0t r=%2d L=%08h R=%08h f=%08h key=%012h",
//                  $time, des_round, des_L, des_R, des_f, des_curkey);
//     end
// end

// // 在 IP 完成那一拍觀察 ip_out, text_in
// always @(posedge clk) begin
//     if (fn_sel == 3'd1 && x == 0 && des_state == 2'd2 && des_round == 0) begin
//         $display("[DES IP] t=%0t text_in=%016h ip_out=%016h",
//                  $time, des_text_in, des_ip_out);
//     end
// end

// `endif
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%



initial begin
   cycle_count = 0;
   @(negedge clk);
   while (1) begin
      cycle_count = cycle_count + 1;
      @(negedge clk);
   end
end


`ifdef p1
   initial begin 
      pattern_file_path = "../00_TESTBED/pattern1_data/pattern1.dat";
      // $display("Hello");
      // $display("%s", pattern_file_path);
      $readmemh(pattern_file_path, pat_mem);
   end
`elsif p2
   initial begin 
      pattern_file_path = "../00_TESTBED/pattern2_data/pattern2.dat";
      $readmemh(pattern_file_path, pat_mem);
   end
`else
   initial begin 
      pattern_file_path = "../00_TESTBED/pattern1_data/pattern1.dat";
      $display("%s", pattern_file_path);
      $readmemh(pattern_file_path, pat_mem);
   end
`endif


`ifdef SDF
   initial       `ifdef SDF_ANNOTATE
   $sdf_annotate(`SDFFILE, u_IOTDF );
`endif
`endif

// initial	 $readmemh("%s/pattern1.dat", pattern_file_path, pat_mem);

`ifdef F2
   initial begin
      func_ans_path = {pattern_file_path[40*8-1:12*8], "f2.dat"};
      $readmemh(func_ans_path, f2_mem); 
      fn_sel=3'd2;  
   end
`elsif F3
   initial begin 
      func_ans_path = {pattern_file_path[40*8-1:12*8], "f3.dat"};
      $readmemh(func_ans_path, f3_mem); 
      fn_sel=3'd3;  
   end
`elsif F4
   initial begin 
      func_ans_path = {pattern_file_path[40*8-1:12*8], "f4.dat"};
      
      $readmemh(func_ans_path, f4_mem); 
      fn_sel=3'd4;  
   end
`else //F1
   initial begin 
      func_ans_path = {pattern_file_path[40*8-1:12*8], "f1.dat"};
      // $display("%s", func_ans_path);
      // $display("%s", pattern_file_path[40*8-1:12*8]);
      $readmemh(func_ans_path, f1_mem); 
      fn_sel=3'd1;  
   end
`endif


initial begin
   clk           = 1'b0;   
   rst           = 1'b0;
   in_en         = 1'b0;   
   i             = 0;
   j             = 15;
   x             = 0;
   in_l          = 0;
   out_h         = 0;
   out_l         = 0;
   pass          = 0;
   err           = 0;
   err_a         = 0;
   over          = 0;
   over1         = 0;
   over2         = 0;
end

always begin #(`CYCLE/2)  clk = ~clk; end

`ifdef vcd
   initial begin
   `ifdef F2
   $dumpfile("IOTDF_F2.vcd");
   `elsif F3
   $dumpfile("IOTDF_F3.vcd");
   `elsif F4
   $dumpfile("IOTDF_F4.vcd");
   `else
   $dumpfile("IOTDF_F1.vcd");
   `endif
   $dumpvars;
   end
`else
   initial begin
   `ifdef F2
   $fsdbDumpfile("IOTDF_F2.fsdb");
   `elsif F3
   $fsdbDumpfile("IOTDF_F3.fsdb");
   `elsif F4
   $fsdbDumpfile("IOTDF_F4.fsdb");
   `else
   $fsdbDumpfile("IOTDF_F1.fsdb");
   `endif
   $fsdbDumpvars;
   $fsdbDumpMDA;
   end
`endif

initial begin
   @(posedge clk)  #`DEL  rst = 1'b1;
   #`CYCLE                rst = 1'b0;

    $display("-----------------------------------------------------\n");  
    $display("Start to Send IOT Data & Compare ...");       
    $display("\n");       
   @(posedge clk)  ;
    while (i < PAT_NUM) begin
      if(!busy)begin     
         in_tmp   = pat_mem[i];
         in_l=127 - j*8; // j is begin from 15

         #`DEL;
         iot_in   =   in_tmp[in_l -: 8];
         // $display("P%02d:  iot_in=%02h, in_tmp[in_l -: 8] =  %02h", x, iot_in, in_tmp[in_l -: 8]);
         in_en    =   1'b1;  

         if(j>0)     j=j-1;
         else begin
                      j=15;
                      i=i+1;              
         end
      end
      else begin
         #`DEL;
         iot_in   = 8'h0;
         in_en    = 1'b0;  
      end
      @(posedge clk);  
    end
    if(busy)begin
	      #`DEL;
         iot_in   = 8'h0;          
    	   in_en    = 1'b0;
    end
    over1 = 1; 
end


always @(posedge clk)begin
   if(valid)begin        
      `ifdef F2
         out_tmp=f2_mem[x];
      `elsif F3
         out_tmp=f3_mem[x];
      `elsif F4
         out_tmp=f4_mem[x];
      `else //F1
         out_tmp=f1_mem[x];
      `endif


      if(iot_out !== out_tmp)begin
         $display("P%02d:  iot_out=%032h  != expect %032h", x, iot_out, out_tmp);
         err = err + 1 ;  
      end
      else begin
         $display("P%02d:  ** Correct!! ** , iot_out=%032h", x, iot_out);
         pass = pass + 1;
      end


         x = x+1;      

      
     `ifdef F2
      if(x >  F2_NUM-1)   over2=1;
     `elsif F3
      if(x >  F3_NUM-1)   over2=1;
     `elsif F4
      if(x >  F4_NUM-1)   over2=1; 
     `else  //F1
      if(x >  F1_NUM-1)   over2=1; 
     `endif

   end                                                                        
end

// // ==== CRC debug：列出 crc_reg 的中間值 ====
// always @(posedge clk) begin
//    // 只在 F3 模式、且 CRC 核心正在跑的時候印
// `ifdef F3
//    if (u_IOTDF.u_crc3_core.running) begin
//       $display("  [CRC dbg] time=%0t  bit_idx=%3d  crc_reg=%03b  data_bit=%b",
//                $time,
//                u_IOTDF.u_crc3_core.bit_idx,
//                u_IOTDF.u_crc3_core.crc_reg,
//                u_IOTDF.u_crc3_core.data_in[u_IOTDF.u_crc3_core.bit_idx]);
//    end
// `endif
// end

always @(*)begin
   over = over1 && over2;
end

initial begin
      @(posedge over)      
      if((over) && (pass !== 'd0) ) begin
         $display("\n-----------------------------------------------------\n");
         if (err == 0)  begin
            $display("Total cost time: %10.2f ns", cycle_count*(`CYCLE));
            
  $display("\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;179;48;5;179m▓\033[38;5;179;48;5;179m▓\033[38;5;173;48;5;173m▓\033[38;5;173;48;5;173m▓\033[38;5;137;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;137;48;5;137m▓\033[38;5;95;48;5;95m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;90;48;5;90m▓\033[38;5;127;48;5;127m▓\033[38;5;91;48;5;91m▓\033[38;5;91;48;5;91m▓\033[38;5;91;48;5;91m▓\033[38;5;127;48;5;127m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;127;48;5;127m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;127;48;5;127m▓\033[38;5;127;48;5;127m▓\033[38;5;91;48;5;91m▓\033[38;5;90;48;5;90m▓\033[38;5;91;48;5;91m▓\033[38;5;90;48;5;90m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;90;48;5;90m▓\033[38;5;132;48;5;132m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;176;48;5;176m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;126;48;5;126m▓\033[0m");
  $display("\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;143;48;5;143m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;179;48;5;179m▓\033[38;5;173;48;5;173m▓\033[38;5;173;48;5;173m▓\033[38;5;137;48;5;137m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;91;48;5;91m▓\033[38;5;127;48;5;127m▓\033[38;5;127;48;5;127m▓\033[38;5;127;48;5;127m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;127;48;5;127m▓\033[38;5;91;48;5;91m▓\033[38;5;91;48;5;91m▓\033[38;5;91;48;5;91m▓\033[38;5;90;48;5;90m▓\033[38;5;90;48;5;90m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;182;48;5;182m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;90;48;5;90m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;126;48;5;126m▓\033[38;5;89;48;5;89m▓\033[0m");
  $display("\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;101;48;5;101m▓\033[38;5;143;48;5;143m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;179;48;5;179m▓\033[38;5;173;48;5;173m▓\033[38;5;137;48;5;137m▓\033[38;5;179;48;5;179m▓\033[38;5;222;48;5;222m▓\033[38;5;186;48;5;186m▓\033[38;5;179;48;5;179m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;90;48;5;90m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;65;48;5;65m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;100;48;5;100m▓\033[38;5;144;48;5;144m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;182;48;5;182m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;53;48;5;53m▓\033[38;5;89;48;5;89m▓\033[38;5;125;48;5;125m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;126;48;5;126m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;143;48;5;143m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;101;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;89;48;5;89m▓\033[38;5;53;48;5;53m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;59;48;5;59m▓\033[38;5;101;48;5;101m▓\033[38;5;137;48;5;137m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;195;48;5;195m▓\033[38;5;231;48;5;231m▓\033[38;5;66;48;5;66m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;109;48;5;109m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;59;48;5;59m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;24;48;5;24m▓\033[38;5;66;48;5;66m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;195;48;5;195m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;95;48;5;95m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;95;48;5;95m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;195;48;5;195m▓\033[38;5;109;48;5;109m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;152;48;5;152m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;126;48;5;126m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;195;48;5;195m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;96;48;5;96m▓\033[38;5;139;48;5;139m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;125;48;5;125m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;125;48;5;125m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;181;48;5;181m▓\033[38;5;96;48;5;96m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;53;48;5;53m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[38;5;126;48;5;126m▓\033[38;5;125;48;5;125m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;109;48;5;109m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;53;48;5;53m▓\033[38;5;125;48;5;125m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;125;48;5;125m▓\033[38;5;125;48;5;125m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;125;48;5;125m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;125;48;5;125m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;168;48;5;168m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;146;48;5;146m▓\033[38;5;67;48;5;67m▓\033[38;5;103;48;5;103m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;53;48;5;53m▓\033[38;5;53;48;5;53m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;139;48;5;139m▓\033[38;5;67;48;5;67m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;60;48;5;60m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;96;48;5;96m▓\033[38;5;132;48;5;132m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;188;48;5;188m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;131;48;5;131m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;53;48;5;53m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;103;48;5;103m▓\033[38;5;146;48;5;146m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;225;48;5;225m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;53;48;5;53m▓\033[38;5;59;48;5;59m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;53;48;5;53m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;110;48;5;110m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;224;48;5;224m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;67;48;5;67m▓\033[38;5;24;48;5;24m▓\033[38;5;17;48;5;17m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;138;48;5;138m▓\033[38;5;59;48;5;59m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;66;48;5;66m▓\033[38;5;67;48;5;67m▓\033[38;5;24;48;5;24m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;67;48;5;67m▓\033[38;5;67;48;5;67m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;96;48;5;96m▓\033[38;5;145;48;5;145m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;96;48;5;96m▓\033[38;5;18;48;5;18m▓\033[38;5;67;48;5;67m▓\033[38;5;24;48;5;24m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;97;48;5;97m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;59;48;5;59m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;67;48;5;67m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;24;48;5;24m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;188;48;5;188m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;96;48;5;96m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;67;48;5;67m▓\033[38;5;60;48;5;60m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;24;48;5;24m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;139;48;5;139m▓\033[38;5;53;48;5;53m▓\033[38;5;133;48;5;133m▓\033[38;5;96;48;5;96m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;132;48;5;132m▓\033[38;5;96;48;5;96m▓\033[38;5;133;48;5;133m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;139;48;5;139m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;67;48;5;67m▓\033[38;5;66;48;5;66m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;139;48;5;139m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;225;48;5;225m▓\033[38;5;181;48;5;181m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;60;48;5;60m▓\033[38;5;24;48;5;24m▓\033[38;5;67;48;5;67m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;96;48;5;96m▓\033[38;5;146;48;5;146m▓\033[38;5;225;48;5;225m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;30;48;5;30m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;53;48;5;53m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;175;48;5;175m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;133;48;5;133m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;97;48;5;97m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;182;48;5;182m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;73;48;5;73m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;96;48;5;96m▓\033[38;5;225;48;5;225m▓\033[38;5;103;48;5;103m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;132;48;5;132m▓\033[38;5;139;48;5;139m▓\033[38;5;138;48;5;138m▓\033[38;5;132;48;5;132m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;54;48;5;54m▓\033[38;5;182;48;5;182m▓\033[38;5;102;48;5;102m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;139;48;5;139m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;132;48;5;132m▓\033[38;5;139;48;5;139m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;60;48;5;60m▓\033[38;5;181;48;5;181m▓\033[38;5;132;48;5;132m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;143;48;5;143m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;142;48;5;142m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;218;48;5;218m▓\033[38;5;54;48;5;54m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;53;48;5;53m▓\033[38;5;89;48;5;89m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;149;48;5;149m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;54;48;5;54m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;139;48;5;139m▓\033[38;5;78;48;5;78m▓\033[38;5;79;48;5;79m▓\033[38;5;67;48;5;67m▓\033[38;5;24;48;5;24m▓\033[38;5;24;48;5;24m▓\033[38;5;67;48;5;67m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;95;48;5;95m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;181;48;5;181m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;182;48;5;182m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;142;48;5;142m▓\033[38;5;142;48;5;142m▓\033[38;5;100;48;5;100m▓\033[38;5;58;48;5;58m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;188;48;5;188m▓\033[38;5;217;48;5;217m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;138;48;5;138m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;189;48;5;189m▓\033[38;5;181;48;5;181m▓\033[38;5;59;48;5;59m▓\033[38;5;115;48;5;115m▓\033[38;5;231;48;5;231m▓\033[38;5;194;48;5;194m▓\033[38;5;157;48;5;157m▓\033[38;5;79;48;5;79m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;60;48;5;60m▓\033[38;5;53;48;5;53m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;182;48;5;182m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;53;48;5;53m▓\033[38;5;103;48;5;103m▓\033[38;5;97;48;5;97m▓\033[38;5;55;48;5;55m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;97;48;5;97m▓\033[38;5;183;48;5;183m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;66;48;5;66m▓\033[38;5;138;48;5;138m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;53;48;5;53m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;53;48;5;53m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;175;48;5;175m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;231;48;5;231m▓\033[38;5;132;48;5;132m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;218;48;5;218m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;188;48;5;188m▓\033[38;5;189;48;5;189m▓\033[38;5;182;48;5;182m▓\033[38;5;140;48;5;140m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;138;48;5;138m▓\033[38;5;224;48;5;224m▓\033[38;5;139;48;5;139m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;188;48;5;188m▓\033[38;5;175;48;5;175m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;140;48;5;140m▓\033[38;5;146;48;5;146m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;224;48;5;224m▓\033[38;5;54;48;5;54m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;132;48;5;132m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;140;48;5;140m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;132;48;5;132m▓\033[38;5;53;48;5;53m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;54;48;5;54m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;60;48;5;60m▓\033[38;5;53;48;5;53m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;89;48;5;89m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;139;48;5;139m▓\033[38;5;61;48;5;61m▓\033[38;5;60;48;5;60m▓\033[38;5;103;48;5;103m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;53;48;5;53m▓\033[38;5;139;48;5;139m▓\033[38;5;132;48;5;132m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;97;48;5;97m▓\033[38;5;146;48;5;146m▓\033[38;5;225;48;5;225m▓\033[38;5;96;48;5;96m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;146;48;5;146m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;89;48;5;89m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;53;48;5;53m▓\033[38;5;96;48;5;96m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;146;48;5;146m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;182;48;5;182m▓\033[38;5;96;48;5;96m▓\033[38;5;97;48;5;97m▓\033[38;5;103;48;5;103m▓\033[38;5;146;48;5;146m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;183;48;5;183m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;53;48;5;53m▓\033[38;5;53;48;5;53m▓\033[38;5;16;48;5;16m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;174;48;5;174m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;102;48;5;102m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;103;48;5;103m▓\033[38;5;97;48;5;97m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;60;48;5;60m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;217;48;5;217m▓\033[38;5;132;48;5;132m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;146;48;5;146m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;61;48;5;61m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;97;48;5;97m▓\033[38;5;225;48;5;225m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;29;48;5;29m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;54;48;5;54m▓\033[38;5;104;48;5;104m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;140;48;5;140m▓\033[38;5;140;48;5;140m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;53;48;5;53m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;29;48;5;29m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;133;48;5;133m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;146;48;5;146m▓\033[38;5;60;48;5;60m▓\033[38;5;189;48;5;189m▓\033[38;5;224;48;5;224m▓\033[38;5;103;48;5;103m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;225;48;5;225m▓\033[38;5;97;48;5;97m▓\033[38;5;145;48;5;145m▓\033[38;5;140;48;5;140m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;132;48;5;132m▓\033[38;5;139;48;5;139m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;139;48;5;139m▓\033[38;5;54;48;5;54m▓\033[38;5;53;48;5;53m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;103;48;5;103m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;183;48;5;183m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;146;48;5;146m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;133;48;5;133m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;95;48;5;95m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;103;48;5;103m▓\033[38;5;183;48;5;183m▓\033[38;5;225;48;5;225m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;61;48;5;61m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;61;48;5;61m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;146;48;5;146m▓\033[38;5;183;48;5;183m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;97;48;5;97m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;72;48;5;72m▓\033[38;5;66;48;5;66m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;98;48;5;98m▓\033[38;5;189;48;5;189m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;97;48;5;97m▓\033[38;5;140;48;5;140m▓\033[38;5;97;48;5;97m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;97;48;5;97m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;96;48;5;96m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;66;48;5;66m▓\033[38;5;72;48;5;72m▓\033[38;5;65;48;5;65m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;97;48;5;97m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;139;48;5;139m▓\033[38;5;61;48;5;61m▓\033[38;5;103;48;5;103m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;59;48;5;59m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;180;48;5;180m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;29;48;5;29m▓\033[38;5;72;48;5;72m▓\033[38;5;66;48;5;66m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;140;48;5;140m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;97;48;5;97m▓\033[38;5;103;48;5;103m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;103;48;5;103m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;60;48;5;60m▓\033[38;5;103;48;5;103m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;103;48;5;103m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;60;48;5;60m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;66;48;5;66m▓\033[38;5;72;48;5;72m▓\033[38;5;72;48;5;72m▓\033[38;5;66;48;5;66m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;140;48;5;140m▓\033[38;5;97;48;5;97m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;139;48;5;139m▓\033[38;5;61;48;5;61m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;53;48;5;53m▓\033[38;5;146;48;5;146m▓\033[38;5;188;48;5;188m▓\033[38;5;139;48;5;139m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;100;48;5;100m▓\033[38;5;100;48;5;100m▓\033[38;5;100;48;5;100m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;217;48;5;217m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;59;48;5;59m▓\033[38;5;72;48;5;72m▓\033[38;5;72;48;5;72m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;96;48;5;96m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;103;48;5;103m▓\033[38;5;140;48;5;140m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;97;48;5;97m▓\033[38;5;61;48;5;61m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;53;48;5;53m▓\033[38;5;60;48;5;60m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;58;48;5;58m▓\033[38;5;142;48;5;142m▓\033[38;5;149;48;5;149m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;143;48;5;143m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;108;48;5;108m▓\033[38;5;66;48;5;66m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;189;48;5;189m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;96;48;5;96m▓\033[38;5;61;48;5;61m▓\033[38;5;104;48;5;104m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;96;48;5;96m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;100;48;5;100m▓\033[38;5;64;48;5;64m▓\033[38;5;64;48;5;64m▓\033[38;5;185;48;5;185m▓\033[38;5;64;48;5;64m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;60;48;5;60m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;60;48;5;60m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;176;48;5;176m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;55;48;5;55m▓\033[38;5;55;48;5;55m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;152;48;5;152m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;146;48;5;146m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;108;48;5;108m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;104;48;5;104m▓\033[38;5;189;48;5;189m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;151;48;5;151m▓\033[38;5;108;48;5;108m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;174;48;5;174m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;60;48;5;60m▓\033[38;5;24;48;5;24m▓\033[38;5;61;48;5;61m▓\033[38;5;67;48;5;67m▓\033[38;5;146;48;5;146m▓\033[38;5;146;48;5;146m▓\033[38;5;189;48;5;189m▓\033[38;5;195;48;5;195m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;97;48;5;97m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;145;48;5;145m▓\033[38;5;108;48;5;108m▓\033[38;5;72;48;5;72m▓\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;59;48;5;59m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;54;48;5;54m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;53;48;5;53m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;72;48;5;72m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;72;48;5;72m▓\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;60;48;5;60m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;103;48;5;103m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;175;48;5;175m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;175;48;5;175m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;139;48;5;139m▓\033[38;5;181;48;5;181m▓\033[38;5;189;48;5;189m▓\033[38;5;146;48;5;146m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;60;48;5;60m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;53;48;5;53m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;139;48;5;139m▓\033[38;5;96;48;5;96m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;61;48;5;61m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;54;48;5;54m▓\033[38;5;18;48;5;18m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;53;48;5;53m▓\033[38;5;132;48;5;132m▓\033[38;5;132;48;5;132m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;188;48;5;188m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;17;48;5;17m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;189;48;5;189m▓\033[38;5;146;48;5;146m▓\033[38;5;103;48;5;103m▓\033[38;5;146;48;5;146m▓\033[38;5;181;48;5;181m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;58;48;5;58m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;131;48;5;131m▓\033[38;5;96;48;5;96m▓\033[38;5;138;48;5;138m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;185;48;5;185m▓\033[38;5;100;48;5;100m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;109;48;5;109m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;175;48;5;175m▓\033[38;5;96;48;5;96m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;136;48;5;136m▓\033[38;5;179;48;5;179m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;221;48;5;221m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;221;48;5;221m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;109;48;5;109m▓\033[38;5;195;48;5;195m▓\033[38;5;195;48;5;195m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;139;48;5;139m▓\033[38;5;133;48;5;133m▓\033[38;5;133;48;5;133m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;132;48;5;132m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;94m▓\033[38;5;179;48;5;179m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;229;48;5;229m▓\033[38;5;185;48;5;185m▓\033[38;5;221;48;5;221m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;136;48;5;136m▓\033[38;5;136;48;5;136m▓\033[38;5;178;48;5;178m▓\033[38;5;221;48;5;221m▓\033[38;5;221;48;5;221m▓\033[38;5;221;48;5;221m▓\033[38;5;100;48;5;100m▓\033[38;5;58;48;5;58m▓\033[38;5;94;48;5;94m▓\033[38;5;100;48;5;100m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;231;48;5;231m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;175;48;5;175m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;139;48;5;139m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;97;48;5;97m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;131;48;5;131m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;229;48;5;229m▓\033[38;5;222;48;5;222m▓\033[38;5;215;48;5;215m▓\033[38;5;221;48;5;221m▓\033[38;5;222;48;5;222m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;222;48;5;222m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;222;48;5;222m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;221;48;5;221m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;179;48;5;179m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;221;48;5;221m▓\033[38;5;58;48;5;58m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;175;48;5;175m▓\033[38;5;133;48;5;133m▓\033[38;5;139;48;5;139m▓\033[38;5;225;48;5;225m▓\033[38;5;175;48;5;175m▓\033[38;5;139;48;5;139m▓\033[38;5;146;48;5;146m▓\033[38;5;224;48;5;224m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;218;48;5;218m▓\033[38;5;183;48;5;183m▓\033[38;5;218;48;5;218m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;216;48;5;216m▓\033[38;5;222;48;5;222m▓\033[38;5;222;48;5;222m▓\033[38;5;216;48;5;216m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;175;48;5;175m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;175;48;5;175m▓\033[38;5;180;48;5;180m▓\033[38;5;221;48;5;221m▓\033[38;5;221;48;5;221m▓\033[38;5;228;48;5;228m▓\033[38;5;222;48;5;222m▓\033[38;5;216;48;5;216m▓\033[38;5;215;48;5;215m▓\033[38;5;179;48;5;179m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;209;48;5;209m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;228;48;5;228m▓\033[38;5;185;48;5;185m▓\033[38;5;172;48;5;172m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;173;48;5;173m▓\033[38;5;173;48;5;173m▓\033[38;5;215;48;5;215m▓\033[38;5;179;48;5;179m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;221;48;5;221m▓\033[38;5;100;48;5;100m▓\033[38;5;58;48;5;58m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;182;48;5;182m▓\033[38;5;133;48;5;133m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;182;48;5;182m▓\033[38;5;139;48;5;139m▓\033[38;5;231;48;5;231m▓\033[38;5;183;48;5;183m▓\033[38;5;133;48;5;133m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;189;48;5;189m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;217;48;5;217m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;179;48;5;179m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;209;48;5;209m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;221;48;5;221m▓\033[38;5;221;48;5;221m▓\033[38;5;228;48;5;228m▓\033[38;5;221;48;5;221m▓\033[38;5;185;48;5;185m▓\033[38;5;179;48;5;179m▓\033[38;5;172;48;5;172m▓\033[38;5;173;48;5;173m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;178;48;5;178m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;221;48;5;221m▓\033[38;5;221;48;5;221m▓\033[38;5;221;48;5;221m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;66;48;5;66m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;181;48;5;181m▓\033[38;5;175;48;5;175m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;218;48;5;218m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;225;48;5;225m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;225;48;5;225m▓\033[38;5;176;48;5;176m▓\033[38;5;225;48;5;225m▓\033[38;5;176;48;5;176m▓\033[38;5;189;48;5;189m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;225;48;5;225m▓\033[38;5;189;48;5;189m▓\033[38;5;189;48;5;189m▓\033[38;5;140;48;5;140m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;140;48;5;140m▓\033[38;5;225;48;5;225m▓\033[38;5;183;48;5;183m▓\033[38;5;225;48;5;225m▓\033[38;5;183;48;5;183m▓\033[38;5;140;48;5;140m▓\033[38;5;139;48;5;139m▓\033[38;5;182;48;5;182m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;218;48;5;218m▓\033[38;5;216;48;5;216m▓\033[38;5;228;48;5;228m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;221;48;5;221m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;222;48;5;222m▓\033[38;5;215;48;5;215m▓\033[38;5;172;48;5;172m▓\033[38;5;221;48;5;221m▓\033[38;5;222;48;5;222m▓\033[38;5;222;48;5;222m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;221;48;5;221m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;228;48;5;228m▓\033[38;5;222;48;5;222m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;215;48;5;215m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;228;48;5;228m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;132;48;5;132m▓\033[38;5;131;48;5;131m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;179;48;5;179m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;185;48;5;185m▓\033[38;5;142;48;5;142m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;22;48;5;22m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;66;48;5;66m▓\033[38;5;29;48;5;29m▓\033[0m");
                  end
         else begin
            $display("Final Simulation Result as below: \n");         
            $display("-----------------------------------------------------\n");
            $display("Pass:   %3d \n", pass);
            $display("Error:  %3d \n", err);
            $display("-----------------------------------------------------\n");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;89;48;5;89m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;94;48;5;94m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;139;48;5;139m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;59;48;5;59m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;109;48;5;109m▓\033[38;5;109;48;5;109m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;167;48;5;167m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;103;48;5;103m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;137;48;5;137m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;175;48;5;175m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;137;48;5;137m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;173;48;5;173m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;223m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;137;48;5;137m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;173;48;5;173m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;173;48;5;173m▓\033[38;5;173;48;5;173m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;94;48;5;94m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;52;48;5;52m▓\033[38;5;94;48;5;94m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;52;48;5;52m▓\033[38;5;58;48;5;58m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;137;48;5;137m▓\033[38;5;174;48;5;174m▓\033[38;5;173;48;5;173m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;137;48;5;137m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;137;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;223;48;5;223m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;95;48;5;95m▓\033[38;5;180;48;5;180m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;225;48;5;225m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;187;48;5;187m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;173;48;5;173m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;137;48;5;137m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;173;48;5;173m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;137;48;5;137m▓\033[38;5;101;48;5;101m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;102;48;5;102m▓\033[38;5;144;48;5;144m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;101;48;5;101m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;131;48;5;131m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;131;48;5;131m▓\033[38;5;138;48;5;138m▓\033[38;5;59;48;5;59m▓\033[38;5;95;48;5;95m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;175;48;5;175m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;146;48;5;146m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;181;48;5;181m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;187;48;5;187m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;95;48;5;95m▓\033[38;5;58;48;5;58m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;59;48;5;59m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;223;48;5;223m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;101;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;180;48;5;180m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;58;48;5;58m▓\033[38;5;94;48;5;94m▓\033[38;5;52;48;5;52m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;109;48;5;109m▓\033[38;5;109;48;5;109m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;103;48;5;103m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;137;48;5;137m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;58;48;5;58m▓\033[38;5;52;48;5;52m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;52;48;5;52m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;187;48;5;187m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;223;48;5;223m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;52;48;5;52m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;95;48;5;95m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;136;48;5;136m▓\033[38;5;173;48;5;173m▓\033[38;5;222;48;5;222m▓\033[38;5;222;48;5;222m▓\033[38;5;58;48;5;58m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;137;48;5;137m▓\033[38;5;94;48;5;94m▓\033[38;5;94;48;5;94m▓\033[38;5;130;48;5;130m▓\033[38;5;94;48;5;94m▓\033[38;5;130;48;5;130m▓\033[38;5;172;48;5;172m▓\033[38;5;215;48;5;215m▓\033[38;5;222;48;5;222m▓\033[38;5;58;48;5;58m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;137;48;5;137m▓\033[38;5;222;48;5;222m▓\033[38;5;216;48;5;216m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;229;48;5;229m▓\033[38;5;229;48;5;229m▓\033[38;5;186;48;5;186m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;103;48;5;103m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;89;48;5;89m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;125;48;5;125m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;52;48;5;52m▓\033[38;5;180;48;5;180m▓\033[38;5;179;48;5;179m▓\033[38;5;222;48;5;222m▓\033[38;5;223;48;5;223m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;58;48;5;58m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;223m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;58;48;5;58m▓\033[38;5;145;48;5;145m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;58;48;5;58m▓\033[38;5;187;48;5;187m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;124;48;5;124m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;52;48;5;52m▓\033[38;5;180;48;5;180m▓\033[38;5;223;48;5;223m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;58;48;5;58m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;132;48;5;132m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;223;48;5;223m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;94;48;5;94m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;223;48;5;223m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;95;48;5;95m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;130;48;5;130m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;131;48;5;131m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;223m▓\033[38;5;144;48;5;144m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;173;48;5;173m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;124;48;5;124m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;180;48;5;180m▓\033[38;5;223;48;5;223m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;131;48;5;131m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;125;48;5;125m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;174;48;5;174m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;131;48;5;131m▓\033[38;5;95;48;5;95m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;174;48;5;174m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;101;48;5;101m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;173;48;5;173m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;95;48;5;95m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;138;48;5;138m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;173;48;5;173m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;210;48;5;210m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;131;48;5;131m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;137;48;5;137m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;130;48;5;130m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;173;48;5;173m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;137;48;5;137m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;125;48;5;125m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;217;48;5;217m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;125;48;5;125m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;60;48;5;60m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;137;48;5;137m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;180;48;5;180m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;53;48;5;53m▓\033[38;5;96;48;5;96m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;137;48;5;137m▓\033[38;5;216;48;5;216m▓\033[38;5;124;48;5;124m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;223;48;5;223m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;180;48;5;180m▓\033[38;5;94;48;5;94m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;53;48;5;53m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;60;48;5;60m▓\033[0m");
  $display("\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;101;48;5;101m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;124;48;5;124m▓\033[38;5;131;48;5;131m▓\033[38;5;181;48;5;181m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[0m");
  $display("\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;95;48;5;95m▓\033[38;5;180;48;5;180m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;124;48;5;124m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;94;48;5;94m▓\033[38;5;130;48;5;130m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;137;48;5;137m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;53;48;5;53m▓\033[38;5;59;48;5;59m▓\033[38;5;95;48;5;95m▓\033[38;5;59;48;5;59m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;59;48;5;59m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;52;48;5;52m▓\033[38;5;131;48;5;131m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;131;48;5;131m▓\033[38;5;124;48;5;124m▓\033[38;5;216;48;5;216m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;223m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;53;48;5;53m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[0m");
  $display("\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;182;48;5;182m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;146;48;5;146m▓\033[38;5;146;48;5;146m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;167;48;5;167m▓\033[38;5;174;48;5;174m▓\033[38;5;94;48;5;94m▓\033[38;5;88;48;5;88m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;17;48;5;17m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[38;5;23;48;5;23m▓\033[0m");
  $display("\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;59;48;5;59m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;216;48;5;216m▓\033[38;5;217;48;5;217m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;137;48;5;137m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;139;48;5;139m▓\033[38;5;95;48;5;95m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;109;48;5;109m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;109;48;5;109m▓\033[38;5;102;48;5;102m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;109;48;5;109m▓\033[38;5;109;48;5;109m▓\033[38;5;103;48;5;103m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;102;48;5;102m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;130;48;5;130m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;53;48;5;53m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;89;48;5;89m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;59;48;5;59m▓\033[38;5;96;48;5;96m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;145;48;5;145m▓\033[38;5;139;48;5;139m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;216;48;5;216m▓\033[38;5;210;48;5;210m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;146;48;5;146m▓\033[38;5;146;48;5;146m▓\033[38;5;182;48;5;182m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;180;48;5;180m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;137;48;5;137m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;95;48;5;95m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;53;48;5;53m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;180;48;5;180m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;173;48;5;173m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;174;48;5;174m▓\033[38;5;181;48;5;181m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;109;48;5;109m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;145;48;5;145m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;108;48;5;108m▓\033[38;5;151;48;5;151m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;101;48;5;101m▓\033[38;5;180;48;5;180m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;138;48;5;138m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;223;48;5;223m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;109;48;5;109m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;53;48;5;53m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;58;48;5;58m▓\033[38;5;138;48;5;138m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;139;48;5;139m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;186;48;5;186m▓\033[38;5;150;48;5;150m▓\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;108;48;5;108m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;102;48;5;102m▓\033[38;5;94;48;5;94m▓\033[38;5;137;48;5;137m▓\033[38;5;216;48;5;216m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;216;48;5;216m▓\033[38;5;216;48;5;216m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;52;48;5;52m▓\033[38;5;53;48;5;53m▓\033[38;5;102;48;5;102m▓\033[38;5;139;48;5;139m▓\033[38;5;103;48;5;103m▓\033[38;5;103;48;5;103m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;108;48;5;108m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;108;48;5;108m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;107;48;5;107m▓\033[38;5;137;48;5;137m▓\033[38;5;173;48;5;173m▓\033[38;5;174;48;5;174m▓\033[38;5;131;48;5;131m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;58;48;5;58m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;139;48;5;139m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;109;48;5;109m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;108;48;5;108m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;64;48;5;64m▓\033[38;5;101;48;5;101m▓\033[38;5;108;48;5;108m▓\033[38;5;144;48;5;144m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;174;48;5;174m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;108;48;5;108m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;108;48;5;108m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;102;48;5;102m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[0m");
  $display("\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;102;48;5;102m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;138;48;5;138m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;66;48;5;66m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;52m▓\033[38;5;144;48;5;144m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;95;48;5;95m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;100;48;5;100m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;139;48;5;139m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[0m");
  $display("\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;108;48;5;108m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;64;48;5;64m▓\033[38;5;107;48;5;107m▓\033[38;5;150;48;5;150m▓\033[38;5;186;48;5;186m▓\033[38;5;144;48;5;144m▓\033[38;5;101;48;5;101m▓\033[38;5;58;48;5;58m▓\033[38;5;95;48;5;95m▓\033[38;5;137;48;5;137m▓\033[38;5;180;48;5;180m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;95;48;5;95m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;102;48;5;102m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;108;48;5;108m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;180;48;5;180m▓\033[38;5;186;48;5;186m▓\033[0m");
  $display("\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;28;48;5;28m▓\033[38;5;107;48;5;107m▓\033[38;5;186;48;5;186m▓\033[38;5;180;48;5;180m▓\033[38;5;186;48;5;186m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;58;48;5;58m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;130;48;5;130m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;185;48;5;185m▓\033[38;5;143;48;5;143m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;150;48;5;150m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;143;48;5;143m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[0m");
  $display("\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;28;48;5;28m▓\033[38;5;65;48;5;65m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;143;48;5;143m▓\033[38;5;101;48;5;101m▓\033[38;5;64;48;5;64m▓\033[38;5;101;48;5;101m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;131;48;5;131m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;52;48;5;52m▓\033[38;5;88;48;5;88m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;65;48;5;65m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;64;48;5;64m▓\033[38;5;58;48;5;58m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;185;48;5;185m▓\033[0m");
  $display("\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;64;48;5;64m▓\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;28;48;5;28m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;101;48;5;101m▓\033[38;5;64;48;5;64m▓\033[38;5;64;48;5;64m▓\033[38;5;138;48;5;138m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;124;48;5;124m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;95;48;5;95m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;107;48;5;107m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;100;48;5;100m▓\033[0m");
  $display("\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;28;48;5;28m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;64;48;5;64m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;58;48;5;58m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;89;48;5;89m▓\033[38;5;89;48;5;89m▓\033[38;5;88;48;5;88m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;138;48;5;138m▓\033[38;5;145;48;5;145m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;64;48;5;64m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[0m");
  $display("\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;64;48;5;64m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;101;48;5;101m▓\033[38;5;150;48;5;150m▓\033[38;5;150;48;5;150m▓\033[38;5;64;48;5;64m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;58;48;5;58m▓\033[38;5;174;48;5;174m▓\033[38;5;210;48;5;210m▓\033[38;5;173;48;5;173m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;88;48;5;88m▓\033[38;5;95;48;5;95m▓\033[38;5;174;48;5;174m▓\033[38;5;217;48;5;217m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;101;48;5;101m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;138;48;5;138m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;23;48;5;23m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;150;48;5;150m▓\033[38;5;101;48;5;101m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;107;48;5;107m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;143;48;5;143m▓\033[38;5;143;48;5;143m▓\033[38;5;144;48;5;144m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;95;48;5;95m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;174;48;5;174m▓\033[38;5;88;48;5;88m▓\033[38;5;94;48;5;94m▓\033[38;5;95;48;5;95m▓\033[38;5;95;48;5;95m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;145;48;5;145m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;187;48;5;187m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;58;48;5;58m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;101;48;5;101m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;64;48;5;64m▓\033[38;5;58;48;5;58m▓\033[38;5;58;48;5;58m▓\033[38;5;58;48;5;58m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;65;48;5;65m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;187;48;5;187m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;181;48;5;181m▓\033[38;5;180;48;5;180m▓\033[38;5;180;48;5;180m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;187;48;5;187m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;187;48;5;187m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;58;48;5;58m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;65;48;5;65m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;144;48;5;144m▓\033[38;5;107;48;5;107m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;102;48;5;102m▓\033[38;5;151;48;5;151m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;52m▓\033[38;5;145;48;5;145m▓\033[38;5;138;48;5;138m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;58;48;5;58m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;186;48;5;186m▓\033[38;5;186;48;5;186m▓\033[38;5;143;48;5;143m▓\033[38;5;107;48;5;107m▓\033[38;5;107;48;5;107m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;58;48;5;58m▓\033[38;5;145;48;5;145m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;187;48;5;187m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;181;48;5;181m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;230;48;5;230m▓\033[38;5;188;48;5;188m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;102;48;5;102m▓\033[38;5;65;48;5;65m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;58;48;5;58m▓\033[38;5;101;48;5;101m▓\033[38;5;150;48;5;150m▓\033[38;5;150;48;5;150m▓\033[38;5;107;48;5;107m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;64;48;5;64m▓\033[38;5;58;48;5;58m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;64;48;5;64m▓\033[38;5;58;48;5;58m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;102;48;5;102m▓\033[38;5;188;48;5;188m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;187;48;5;187m▓\033[38;5;138;48;5;138m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;194;48;5;194m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;187;48;5;187m▓\033[38;5;144;48;5;144m▓\033[38;5;143;48;5;143m▓\033[38;5;101;48;5;101m▓\033[38;5;65;48;5;65m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;65;48;5;65m▓\033[38;5;65;48;5;65m▓\033[38;5;64;48;5;64m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;65;48;5;65m▓\033[38;5;66;48;5;66m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;145;48;5;145m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;22;48;5;22m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;230;48;5;230m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;144;48;5;144m▓\033[38;5;102;48;5;102m▓\033[38;5;65;48;5;65m▓\033[38;5;22;48;5;22m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;230;48;5;230m▓\033[38;5;188;48;5;188m▓\033[38;5;144;48;5;144m▓\033[38;5;145;48;5;145m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;60;48;5;60m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;60;48;5;60m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;102;48;5;102m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;144;48;5;144m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;102;48;5;102m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;66;48;5;66m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;95;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;101;48;5;101m▓\033[38;5;181;48;5;181m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[0m");
  $display("\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;138;48;5;138m▓\033[38;5;188;48;5;188m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;224;48;5;224m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;181;48;5;181m▓\033[38;5;144;48;5;144m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;138;48;5;138m▓\033[38;5;95;48;5;95m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;60;48;5;60m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;102;48;5;102m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;52m▓\033[38;5;52;48;5;52m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;53;48;5;53m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;65;48;5;65m▓\033[38;5;59;48;5;59m▓\033[38;5;66;48;5;66m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;60;48;5;60m▓\033[38;5;66;48;5;66m▓\033[38;5;66;48;5;66m▓\033[38;5;59;48;5;59m▓\033[38;5;109;48;5;109m▓\033[38;5;151;48;5;151m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;187;48;5;187m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;145;48;5;145m▓\033[38;5;59;48;5;59m▓\033[38;5;59;48;5;59m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;187;48;5;187m▓\033[38;5;181;48;5;181m▓\033[38;5;181;48;5;181m▓\033[0m");
         end
      end
      #(`CYCLE/2); $finish;
end

initial begin
	#(`End_CYCLE*(`CYCLE));
	$display("-----------------------------------------------------\n");
	$display("Error!!! There is something wrong with your code ...!\n");
 	$display("------The test result is .....FAIL ------------------\n");
 	$display("-----------------------------------------------------\n");
 	$finish;
end
   

   
endmodule



