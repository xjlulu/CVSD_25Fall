`timescale 1ns/100ps

module imm_gen (
    input  wire [31:0] i_instr,
    output reg  [31:0] o_imm
);

    wire [6:0] opcode = i_instr[6:0];

    always @(*) begin
        case (opcode)
            // ---------------------------------------------------------------
            // I-type (ADDI, JALR, LW)
            // ---------------------------------------------------------------
            7'b0010011, // ADDI
            7'b1100111, // JALR
            7'b0000111, // FLW
            7'b0000011: // LW
                o_imm = {{20{i_instr[31]}}, i_instr[31:20]}; // sign-extend

            // ---------------------------------------------------------------
            // S-type (SW)
            // ---------------------------------------------------------------
            7'b0100111, // FSW
            7'b0100011:
                o_imm = {{20{i_instr[31]}}, i_instr[31:25], i_instr[11:7]};

            // ---------------------------------------------------------------
            // B-type (BEQ, BLT)
            // ---------------------------------------------------------------
            7'b1100011:
                o_imm = {{20{i_instr[31]}}, i_instr[7],
                         i_instr[30:25], i_instr[11:8], 1'b0};

            // ---------------------------------------------------------------
            // U-type (AUIPC)
            // ---------------------------------------------------------------
            7'b0010111:
                o_imm = {i_instr[31:12], 12'd0};

            // ---------------------------------------------------------------
            // Default: zero immediate
            // ---------------------------------------------------------------
            default:
                o_imm = 32'd0;
        endcase
    end
endmodule
